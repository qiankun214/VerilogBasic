module PLBI2F (
	input CONOF,
	input SONOF,
	input A,
	input E,
	input PU,
	input PD,
	input P,
	input D
);

endmodule