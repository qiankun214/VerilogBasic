
module ROM_4 (
    input [7:0]addr,
    output reg [7:0]dout
);

always @(*) begin
    case(addr)
		8'd0:dout = 8'd0;
		8'd1:dout = 8'd0;
		8'd2:dout = 8'd0;
		8'd3:dout = 8'd0;
		8'd4:dout = 8'd0;
		8'd5:dout = 8'd0;
		8'd6:dout = 8'd0;
		8'd7:dout = 8'd0;
		8'd8:dout = 8'd0;
		8'd9:dout = 8'd0;
		8'd10:dout = 8'd0;
		8'd11:dout = 8'd0;
		8'd12:dout = 8'd0;
		8'd13:dout = 8'd0;
		8'd14:dout = 8'd0;
		8'd15:dout = 8'd0;
		8'd16:dout = 8'd0;
		8'd17:dout = 8'd1;
		8'd18:dout = 8'd2;
		8'd19:dout = 8'd3;
		8'd20:dout = 8'd4;
		8'd21:dout = 8'd5;
		8'd22:dout = 8'd6;
		8'd23:dout = 8'd7;
		8'd24:dout = 8'd8;
		8'd25:dout = 8'd9;
		8'd26:dout = 8'd10;
		8'd27:dout = 8'd11;
		8'd28:dout = 8'd12;
		8'd29:dout = 8'd13;
		8'd30:dout = 8'd14;
		8'd31:dout = 8'd15;
		8'd32:dout = 8'd0;
		8'd33:dout = 8'd2;
		8'd34:dout = 8'd4;
		8'd35:dout = 8'd6;
		8'd36:dout = 8'd8;
		8'd37:dout = 8'd10;
		8'd38:dout = 8'd12;
		8'd39:dout = 8'd14;
		8'd40:dout = 8'd16;
		8'd41:dout = 8'd18;
		8'd42:dout = 8'd20;
		8'd43:dout = 8'd22;
		8'd44:dout = 8'd24;
		8'd45:dout = 8'd26;
		8'd46:dout = 8'd28;
		8'd47:dout = 8'd30;
		8'd48:dout = 8'd0;
		8'd49:dout = 8'd3;
		8'd50:dout = 8'd6;
		8'd51:dout = 8'd9;
		8'd52:dout = 8'd12;
		8'd53:dout = 8'd15;
		8'd54:dout = 8'd18;
		8'd55:dout = 8'd21;
		8'd56:dout = 8'd24;
		8'd57:dout = 8'd27;
		8'd58:dout = 8'd30;
		8'd59:dout = 8'd33;
		8'd60:dout = 8'd36;
		8'd61:dout = 8'd39;
		8'd62:dout = 8'd42;
		8'd63:dout = 8'd45;
		8'd64:dout = 8'd0;
		8'd65:dout = 8'd4;
		8'd66:dout = 8'd8;
		8'd67:dout = 8'd12;
		8'd68:dout = 8'd16;
		8'd69:dout = 8'd20;
		8'd70:dout = 8'd24;
		8'd71:dout = 8'd28;
		8'd72:dout = 8'd32;
		8'd73:dout = 8'd36;
		8'd74:dout = 8'd40;
		8'd75:dout = 8'd44;
		8'd76:dout = 8'd48;
		8'd77:dout = 8'd52;
		8'd78:dout = 8'd56;
		8'd79:dout = 8'd60;
		8'd80:dout = 8'd0;
		8'd81:dout = 8'd5;
		8'd82:dout = 8'd10;
		8'd83:dout = 8'd15;
		8'd84:dout = 8'd20;
		8'd85:dout = 8'd25;
		8'd86:dout = 8'd30;
		8'd87:dout = 8'd35;
		8'd88:dout = 8'd40;
		8'd89:dout = 8'd45;
		8'd90:dout = 8'd50;
		8'd91:dout = 8'd55;
		8'd92:dout = 8'd60;
		8'd93:dout = 8'd65;
		8'd94:dout = 8'd70;
		8'd95:dout = 8'd75;
		8'd96:dout = 8'd0;
		8'd97:dout = 8'd6;
		8'd98:dout = 8'd12;
		8'd99:dout = 8'd18;
		8'd100:dout = 8'd24;
		8'd101:dout = 8'd30;
		8'd102:dout = 8'd36;
		8'd103:dout = 8'd42;
		8'd104:dout = 8'd48;
		8'd105:dout = 8'd54;
		8'd106:dout = 8'd60;
		8'd107:dout = 8'd66;
		8'd108:dout = 8'd72;
		8'd109:dout = 8'd78;
		8'd110:dout = 8'd84;
		8'd111:dout = 8'd90;
		8'd112:dout = 8'd0;
		8'd113:dout = 8'd7;
		8'd114:dout = 8'd14;
		8'd115:dout = 8'd21;
		8'd116:dout = 8'd28;
		8'd117:dout = 8'd35;
		8'd118:dout = 8'd42;
		8'd119:dout = 8'd49;
		8'd120:dout = 8'd56;
		8'd121:dout = 8'd63;
		8'd122:dout = 8'd70;
		8'd123:dout = 8'd77;
		8'd124:dout = 8'd84;
		8'd125:dout = 8'd91;
		8'd126:dout = 8'd98;
		8'd127:dout = 8'd105;
		8'd128:dout = 8'd0;
		8'd129:dout = 8'd8;
		8'd130:dout = 8'd16;
		8'd131:dout = 8'd24;
		8'd132:dout = 8'd32;
		8'd133:dout = 8'd40;
		8'd134:dout = 8'd48;
		8'd135:dout = 8'd56;
		8'd136:dout = 8'd64;
		8'd137:dout = 8'd72;
		8'd138:dout = 8'd80;
		8'd139:dout = 8'd88;
		8'd140:dout = 8'd96;
		8'd141:dout = 8'd104;
		8'd142:dout = 8'd112;
		8'd143:dout = 8'd120;
		8'd144:dout = 8'd0;
		8'd145:dout = 8'd9;
		8'd146:dout = 8'd18;
		8'd147:dout = 8'd27;
		8'd148:dout = 8'd36;
		8'd149:dout = 8'd45;
		8'd150:dout = 8'd54;
		8'd151:dout = 8'd63;
		8'd152:dout = 8'd72;
		8'd153:dout = 8'd81;
		8'd154:dout = 8'd90;
		8'd155:dout = 8'd99;
		8'd156:dout = 8'd108;
		8'd157:dout = 8'd117;
		8'd158:dout = 8'd126;
		8'd159:dout = 8'd135;
		8'd160:dout = 8'd0;
		8'd161:dout = 8'd10;
		8'd162:dout = 8'd20;
		8'd163:dout = 8'd30;
		8'd164:dout = 8'd40;
		8'd165:dout = 8'd50;
		8'd166:dout = 8'd60;
		8'd167:dout = 8'd70;
		8'd168:dout = 8'd80;
		8'd169:dout = 8'd90;
		8'd170:dout = 8'd100;
		8'd171:dout = 8'd110;
		8'd172:dout = 8'd120;
		8'd173:dout = 8'd130;
		8'd174:dout = 8'd140;
		8'd175:dout = 8'd150;
		8'd176:dout = 8'd0;
		8'd177:dout = 8'd11;
		8'd178:dout = 8'd22;
		8'd179:dout = 8'd33;
		8'd180:dout = 8'd44;
		8'd181:dout = 8'd55;
		8'd182:dout = 8'd66;
		8'd183:dout = 8'd77;
		8'd184:dout = 8'd88;
		8'd185:dout = 8'd99;
		8'd186:dout = 8'd110;
		8'd187:dout = 8'd121;
		8'd188:dout = 8'd132;
		8'd189:dout = 8'd143;
		8'd190:dout = 8'd154;
		8'd191:dout = 8'd165;
		8'd192:dout = 8'd0;
		8'd193:dout = 8'd12;
		8'd194:dout = 8'd24;
		8'd195:dout = 8'd36;
		8'd196:dout = 8'd48;
		8'd197:dout = 8'd60;
		8'd198:dout = 8'd72;
		8'd199:dout = 8'd84;
		8'd200:dout = 8'd96;
		8'd201:dout = 8'd108;
		8'd202:dout = 8'd120;
		8'd203:dout = 8'd132;
		8'd204:dout = 8'd144;
		8'd205:dout = 8'd156;
		8'd206:dout = 8'd168;
		8'd207:dout = 8'd180;
		8'd208:dout = 8'd0;
		8'd209:dout = 8'd13;
		8'd210:dout = 8'd26;
		8'd211:dout = 8'd39;
		8'd212:dout = 8'd52;
		8'd213:dout = 8'd65;
		8'd214:dout = 8'd78;
		8'd215:dout = 8'd91;
		8'd216:dout = 8'd104;
		8'd217:dout = 8'd117;
		8'd218:dout = 8'd130;
		8'd219:dout = 8'd143;
		8'd220:dout = 8'd156;
		8'd221:dout = 8'd169;
		8'd222:dout = 8'd182;
		8'd223:dout = 8'd195;
		8'd224:dout = 8'd0;
		8'd225:dout = 8'd14;
		8'd226:dout = 8'd28;
		8'd227:dout = 8'd42;
		8'd228:dout = 8'd56;
		8'd229:dout = 8'd70;
		8'd230:dout = 8'd84;
		8'd231:dout = 8'd98;
		8'd232:dout = 8'd112;
		8'd233:dout = 8'd126;
		8'd234:dout = 8'd140;
		8'd235:dout = 8'd154;
		8'd236:dout = 8'd168;
		8'd237:dout = 8'd182;
		8'd238:dout = 8'd196;
		8'd239:dout = 8'd210;
		8'd240:dout = 8'd0;
		8'd241:dout = 8'd15;
		8'd242:dout = 8'd30;
		8'd243:dout = 8'd45;
		8'd244:dout = 8'd60;
		8'd245:dout = 8'd75;
		8'd246:dout = 8'd90;
		8'd247:dout = 8'd105;
		8'd248:dout = 8'd120;
		8'd249:dout = 8'd135;
		8'd250:dout = 8'd150;
		8'd251:dout = 8'd165;
		8'd252:dout = 8'd180;
		8'd253:dout = 8'd195;
		8'd254:dout = 8'd210;
		8'd255:dout = 8'd225;
		default:dout = 'b0;
    endcase
end
endmodule
